-------------------------------------------------------------------------------
--
-- The IN port controller.
--
-- $Id: t400_io_in-c.vhd,v 1.1 2006-05-22 00:00:55 arniml Exp $
--
-- Copyright (c) 2006, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t400_io_in_rtl_c0 of t400_io_in is

  for rtl
  end for;

end t400_io_in_rtl_c0;


-------------------------------------------------------------------------------
-- File History:
--
-- $Log: not supported by cvs2svn $
-------------------------------------------------------------------------------
