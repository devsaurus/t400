-------------------------------------------------------------------------------
--
-- The serial input/output unit.
--
-- $Id$
--
-- Copyright (c) 2006, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t400_sio_rtl_c0 of t400_sio is

  for rtl
  end for;

end t400_sio_rtl_c0;
