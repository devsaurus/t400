-------------------------------------------------------------------------------
--
-- The Data memory controller.
--
-- $Id$
--
-- Copyright (c) 2006, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t400_dmem_ctrl_rtl_c0 of t400_dmem_ctrl is

  for rtl
  end for;

end t400_dmem_ctrl_rtl_c0;
