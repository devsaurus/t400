-------------------------------------------------------------------------------
--
-- The reset generation unit.
--
-- $Id: t400_reset-c.vhd,v 1.1.1.1 2006-05-06 01:56:45 arniml Exp $
--
-- Copyright (c) 2006, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t400_reset_rtl_c0 of t400_reset is

  for rtl
  end for;

end t400_reset_rtl_c0;


-------------------------------------------------------------------------------
-- File History:
--
-- $Log: not supported by cvs2svn $
-------------------------------------------------------------------------------
