-------------------------------------------------------------------------------
-- $Id: t400_por-c.vhd,v 1.1.1.1 2006-05-06 01:56:44 arniml Exp $
-------------------------------------------------------------------------------

configuration t400_por_cyclone_c0 of t400_por is

  for cyclone
  end for;

end t400_por_cyclone_c0;


-------------------------------------------------------------------------------
-- File History:
--
-- $Log: not supported by cvs2svn $
-------------------------------------------------------------------------------
