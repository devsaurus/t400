-------------------------------------------------------------------------------
--
-- The reset generation unit.
--
-- $Id$
--
-- Copyright (c) 2006, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t400_reset_rtl_c0 of t400_reset is

  for rtl
  end for;

end t400_reset_rtl_c0;
