-------------------------------------------------------------------------------
--
-- Generic testbench elements
--
-- $Id$
--
-- Copyright (c) 2006, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration tb_elems_behav_c0 of tb_elems is

  for behav
  end for;

end tb_elems_behav_c0;
