-------------------------------------------------------------------------------
--
-- The timer unit.
--
-- $Id$
--
-- Copyright (c) 2006, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t400_timer_rtl_c0 of t400_timer is

  for rtl
  end for;

end t400_timer_rtl_c0;
