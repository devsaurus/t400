-------------------------------------------------------------------------------
--
-- The IN port controller.
--
-- $Id$
--
-- Copyright (c) 2006, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t400_io_in_rtl_c0 of t400_io_in is

  for rtl
  end for;

end t400_io_in_rtl_c0;
