-------------------------------------------------------------------------------
-- $Id: t400_por-c.vhd,v 1.1 2006-05-07 01:47:51 arniml Exp $
-------------------------------------------------------------------------------

configuration t400_por_rtl_c0 of t400_por is

  for spartan
  end for;

end t400_por_rtl_c0;


-------------------------------------------------------------------------------
-- File History:
--
-- $Log: not supported by cvs2svn $
-------------------------------------------------------------------------------
