-------------------------------------------------------------------------------
--
-- Generic testbench elements
--
-- $Id: tb_elems-c.vhd,v 1.1 2006-05-15 21:55:27 arniml Exp $
--
-- Copyright (c) 2006, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration tb_elems_behav_c0 of tb_elems is

  for behav
  end for;

end tb_elems_behav_c0;


-------------------------------------------------------------------------------
-- File History:
--
-- $Log: not supported by cvs2svn $
-------------------------------------------------------------------------------
