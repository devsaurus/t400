-------------------------------------------------------------------------------
-- $Id$
-------------------------------------------------------------------------------

configuration t400_por_rtl_c0 of t400_por is

  for cyclone
  end for;

end t400_por_rtl_c0;
