-------------------------------------------------------------------------------
--
-- The L port controller.
--
-- $Id: t400_io_l-c.vhd,v 1.1.1.1 2006-05-06 01:56:44 arniml Exp $
--
-- Copyright (c) 2006, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t400_io_l_rtl_c0 of t400_io_l is

  for rtl
  end for;

end t400_io_l_rtl_c0;


-------------------------------------------------------------------------------
-- File History:
--
-- $Log: not supported by cvs2svn $
-------------------------------------------------------------------------------
