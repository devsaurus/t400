-------------------------------------------------------------------------------
--
-- The timer unit.
--
-- $Id: t400_timer-c.vhd,v 1.1 2006-05-20 02:47:12 arniml Exp $
--
-- Copyright (c) 2006, Arnim Laeuger (arniml@opencores.org)
--
-- All rights reserved
--
-------------------------------------------------------------------------------

configuration t400_timer_rtl_c0 of t400_timer is

  for rtl
  end for;

end t400_timer_rtl_c0;


-------------------------------------------------------------------------------
-- File History:
--
-- $Log: not supported by cvs2svn $
-------------------------------------------------------------------------------
